module uart_tx(
input	logic			clk,
input 	logic			rst_,
input	logic			tx_start,
input	logic	[7:0]	tx_data,
output	logic			tx_serial,
output	logic			tx_busy
);




endmodule 